// Write a verilog code to print hello world
module Second;
initial
    begin
        $display("Hello, World");
        $finish ;
    end
endmodule